module display (
    
    ports
);
    
endmodule