module Debounce(
    input num,
    input clk,
    output num_o, digit
);

    wire clk_div;
    wire q1, q2, nq2, q0;
    wire num;

    FrecDivider ClkDiv(clk, clk_div);

    D_FF KB_i (clk, clk_div, num, q0);
    D_FF KB_FF1(clk, clk_div, q0, q1);
    D_FF KB_FF1(clk, clk_div, q1, q2);

    assign nq2 = ~q2;
    assign num_o = q1 & nq2;
    
    always @(posedge clk_div) begin
        if (num_o = q1 & nq2) begin
            digit = q2;
        end
    end

endmodule